// Defines for ULX3S